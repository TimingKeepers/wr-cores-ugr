library ieee;
use ieee.std_logic_1164.all;


package wr_fabric_pkg is

  constant c_WRF_DATA   : std_logic_vector(1 downto 0) := "00";
  constant c_WRF_OOB    : std_logic_vector(1 downto 0) := "01";
  constant c_WRF_STATUS : std_logic_vector(1 downto 0) := "10";
  constant c_WRF_USER   : std_logic_vector(1 downto 0) := "11";

  constant c_WRF_OOB_TYPE_RX : std_logic_vector(3 downto 0) := "0000";
  constant c_WRF_OOB_TYPE_TX : std_logic_vector(3 downto 0) := "0001";

  type t_wrf_oob is record
    ts_r: std_logic_vector(27 downto 0);
    ts_f: std_logic_vector(3 downto 0);
    port_id: std_logic_vector(5 downto 0);
    frame_id: std_logic_vector(15 downto 0);
  end record;
  
  type t_wrf_status_reg is record
    is_hp       : std_logic;
    has_smac    : std_logic;
    has_crc     : std_logic;
    rx_error    : std_logic;
    tag_me      : std_logic;
    match_class : std_logic_vector(7 downto 0);
  end record;

  type t_wrf_source_out is record
    adr : std_logic_vector(1 downto 0);
    dat : std_logic_vector(15 downto 0);
    cyc : std_logic;
    stb : std_logic;
    we  : std_logic;
    sel : std_logic_vector(1 downto 0);
  end record;

  type t_wrf_source_in is record
    ack   : std_logic;
    stall : std_logic;
  end record;

  subtype t_wrf_sink_in is t_wrf_source_out;
  subtype t_wrf_sink_out is t_wrf_source_in;

  
  function f_marshall_wrf_status (stat  : t_wrf_status_reg) return std_logic_vector;
  function f_unmarshall_wrf_status(stat : std_logic_vector) return t_wrf_status_reg;

  
end wr_fabric_pkg;

package body wr_fabric_pkg is

    function f_marshall_wrf_status(stat : t_wrf_status_reg)
    return std_logic_vector is
    variable tmp : std_logic_vector(15 downto 0);
  begin
    tmp(0)           := stat.is_hp;
    tmp(1)           := stat.rx_error;
    tmp(2)           := stat.has_smac;
    tmp(15 downto 8) := stat.match_class;
    return tmp;
  end function;

  function f_unmarshall_wrf_status(stat : std_logic_vector) return t_wrf_status_reg is
    variable tmp : t_wrf_status_reg;
  begin
    tmp.is_hp       := stat(0);
    tmp.rx_error    := stat(1);
    tmp.has_smac    := stat(2);
    tmp.match_class := stat(15 downto 8);
    return tmp;
    
  end function;


end wr_fabric_pkg;
