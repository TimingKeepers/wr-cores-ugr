dmtd_clk_pll_inst : dmtd_clk_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
