-------------------------------------------------------------------------------
-- Title      : Mini Embedded DMA Network Interface Controller
-- Project    : WhiteRabbit Core
-------------------------------------------------------------------------------
-- File       : wrsw_mini_nic.vhd
-- Author     : Tomasz Wlostowski
-- Company    : CERN BE-Co-HT
-- Created    : 2010-07-26
-- Last update: 2011-10-24
-- Platform   : FPGA-generic
-- Standard   : VHDL
-------------------------------------------------------------------------------
-- Description: Module implements a simple NIC with DMA controller. It
-- sends/receives the packets using WR switch fabric interface (see the
-- wrsw_endpoint.vhd for the details). Packets are stored and read from the
-- system memory via simple memory bus. WR endpoint-compatible TX timestamping
-- unit is also included.
-------------------------------------------------------------------------------
-- Copyright (c) 2010, 2011 CERN
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2010-07-26  1.0      twlostow        Created
-- 2010-08-16  1.0      twlostow        Bugfixes, linux compatibility added
-- 2011-08-03  2.0      greg.d          rewritten to use pipelined Wishbone
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.wr_fabric_pkg.all;
use work.wishbone_pkg.all;
use work.minic_wbgen2_pkg.all;


entity wr_mini_nic is

  generic (
    g_interface_mode       : t_wishbone_interface_mode      := CLASSIC;
    g_address_granularity  : t_wishbone_address_granularity := WORD;
    g_memsize_log2         : integer                        := 14;
    g_buffer_little_endian : boolean                        := true);

  port (
    clk_sys_i : in std_logic;
    rst_n_i   : in std_logic;

-------------------------------------------------------------------------------
-- System memory i/f
-------------------------------------------------------------------------------

    mem_data_o : out std_logic_vector(31 downto 0);
    mem_addr_o : out std_logic_vector(g_memsize_log2-1 downto 0);
    mem_data_i : in  std_logic_vector(31 downto 0);
    mem_wr_o   : out std_logic;

-------------------------------------------------------------------------------
-- Pipelined Wishbone interface
-------------------------------------------------------------------------------

    -- WBP Master (TX)
    src_dat_o   : out std_logic_vector(15 downto 0);
    src_adr_o   : out std_logic_vector(1 downto 0);
    src_sel_o   : out std_logic_vector(1 downto 0);
    src_cyc_o   : out std_logic;
    src_stb_o   : out std_logic;
    src_we_o    : out std_logic;
    src_stall_i : in  std_logic;
    src_err_i   : in  std_logic;
    src_ack_i   : in  std_logic;

    -- WBP Slave (RX)
    snk_dat_i   : in  std_logic_vector(15 downto 0);
    snk_adr_i   : in  std_logic_vector(1 downto 0);
    snk_sel_i   : in  std_logic_vector(1 downto 0);
    snk_cyc_i   : in  std_logic;
    snk_stb_i   : in  std_logic;
    snk_we_i    : in  std_logic;
    snk_stall_o : out std_logic;
    snk_err_o   : out std_logic;
    snk_ack_o   : out std_logic;

-------------------------------------------------------------------------------
-- TXTSU i/f
-------------------------------------------------------------------------------

    txtsu_port_id_i  : in  std_logic_vector(4 downto 0);
    txtsu_frame_id_i : in  std_logic_vector(16 - 1 downto 0);
    txtsu_tsval_i    : in  std_logic_vector(28 + 4 - 1 downto 0);
    txtsu_valid_i    : in  std_logic;
    txtsu_ack_o      : out std_logic;

-------------------------------------------------------------------------------
-- Wishbone slave
-------------------------------------------------------------------------------    

    wb_cyc_i   : in  std_logic;
    wb_stb_i   : in  std_logic;
    wb_we_i    : in  std_logic;
    wb_sel_i   : in  std_logic_vector(c_wishbone_data_width/8-1 downto 0);
    wb_adr_i   : in  std_logic_vector(c_wishbone_address_width-1 downto 0);
    wb_dat_i   : in  std_logic_vector(c_wishbone_data_width-1 downto 0);
    wb_dat_o   : out std_logic_vector(c_wishbone_data_width-1 downto 0);
    wb_ack_o   : out std_logic;
    wb_stall_o : out std_logic;
    wb_irq_o   : out std_logic
    );
end wr_mini_nic;

architecture behavioral of wr_mini_nic is

  component minic_wb_slave
    port (
      rst_n_i          : in  std_logic;
      wb_clk_i         : in  std_logic;
      wb_addr_i        : in  std_logic_vector(3 downto 0);
      wb_data_i        : in  std_logic_vector(31 downto 0);
      wb_data_o        : out std_logic_vector(31 downto 0);
      wb_cyc_i         : in  std_logic;
      wb_sel_i         : in  std_logic_vector(3 downto 0);
      wb_stb_i         : in  std_logic;
      wb_we_i          : in  std_logic;
      wb_ack_o         : out std_logic;
      wb_irq_o         : out std_logic;
      tx_ts_read_ack_o : out std_logic;
      irq_tx_i         : in  std_logic;
      irq_tx_ack_o     : out std_logic;
      irq_tx_mask_o    : out std_logic;
      irq_rx_i         : in  std_logic;
      irq_rx_ack_o     : out std_logic;
      irq_txts_i       : in  std_logic;
      regs_i           : in  t_minic_in_registers;
      regs_o           : out t_minic_out_registers);
  end component;

  type t_wrf_status_reg is record
    is_hp       : std_logic;
    has_smac    : std_logic;
    has_crc     : std_logic;
    error       : std_logic;
    tag_me      : std_logic;
    match_class : std_logic_vector(7 downto 0);
  end record;

  function f_buf_swap_endian_32
    (
      data : std_logic_vector(31 downto 0)
      ) return std_logic_vector is
  begin
    if(g_buffer_little_endian = true) then
      return data(7 downto 0) & data(15 downto 8) & data(23 downto 16) & data(31 downto 24);
    else
      return data;
    end if;
  end function f_buf_swap_endian_32;


-----------------------------------------------------------------------------
-- memory interface signals
-----------------------------------------------------------------------------

  signal ntx_mem_d  : std_logic_vector(31 downto 0);
  signal ntx_mem_a  : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_mem_d  : std_logic_vector(31 downto 0);
  signal nrx_mux_d  : std_logic;
  signal nrx_mem_a  : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_mem_wr : std_logic;
  signal mem_arb_rx : std_logic;
  signal mem_arb_tx : std_logic;


-------------------------------------------------------------------------------
-- TX FSM stuff
-------------------------------------------------------------------------------

  type t_tx_fsm_state is (TX_IDLE, TX_READ_DESC, TX_STATUS, TX_START_PACKET, TX_HWORD, TX_LWORD, TX_END_PACKET);

  alias ntx_desc_size is ntx_mem_d(g_memsize_log2 downto 0);
  alias ntx_desc_odd is ntx_mem_d(0);
  alias ntx_desc_valid is ntx_mem_d(31);
  alias ntx_desc_with_oob is ntx_mem_d(30);
  alias ntx_desc_802_1q is ntx_mem_d(29);
  alias ntx_desc_has_src_mac is ntx_mem_d(28);

  --STATUS Reg for TX path
  signal ntx_status_reg : std_logic_vector(15 downto 0);
  alias ntx_status_class is ntx_status_reg(7 downto 0);
  alias ntx_status_tagme is ntx_status_reg(8);
  alias ntx_status_err is ntx_status_reg(9);
  alias ntx_status_crc is ntx_status_reg(10);
  alias ntx_status_smac is ntx_status_reg(11);
  alias ntx_status_hp is ntx_status_reg(12);

  signal ntx_data_reg : std_logic_vector(31 downto 0);

  signal ntx_cntr_is_zero    : std_logic;
  signal ntx_cntr_is_one     : std_logic;
  signal ntx_ackcntr_is_zero : std_logic;
  signal ntx_timeout_is_zero : std_logic;
  signal ntx_cntr            : unsigned(g_memsize_log2 downto 0);
  signal ntx_ackcntr         : unsigned(g_memsize_log2 downto 0);
  signal ntx_timeout         : unsigned(7 downto 0);
  signal ntx_has_oob         : std_logic;
  signal ntx_state           : t_tx_fsm_state;
  signal ntx_curst           : t_tx_fsm_state;
  signal ntx_start_delayed   : std_logic;
  signal ntx_size_odd        : std_logic;

-------------------------------------------------------------------------------
-- RX FSM stuff
-------------------------------------------------------------------------------  

  type t_rx_fsm_state is (RX_WAIT_SOF, RX_MEM_RESYNC, RX_MEM_FLUSH, RX_ALLOCATE_DESCRIPTOR, RX_DATA, RX_UPDATE_DESC);

  signal nrx_state   : t_rx_fsm_state;
  signal nrx_avail   : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_toggle  : std_logic;
  signal nrx_oob_reg : std_logic_vector(15 downto 0);

  --STATUS Reg for RX path
  signal nrx_status_reg : std_logic_vector(15 downto 0);
  alias nrx_status_class is nrx_status_reg(7 downto 0);
  alias nrx_status_tagme is nrx_status_reg(8);
  alias nrx_status_err is nrx_status_reg(9);
  alias nrx_status_crc is nrx_status_reg(10);
  alias nrx_status_smac is nrx_status_reg(11);
  alias nrx_status_hp is nrx_status_reg(12);

  signal nrx_mem_a_saved : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_has_oob     : std_logic;
  signal nrx_bytesel     : std_logic;
  signal nrx_size        : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_acksize     : unsigned(g_memsize_log2-1 downto 0);
  signal nrx_buf_full    : std_logic;
  signal nrx_stall_mask  : std_logic;

-------------------------------------------------------------------------------
-- Classic Wishbone slave signals
-------------------------------------------------------------------------------  

  signal regs_in  : t_minic_in_registers;
  signal regs_out : t_minic_out_registers;

  signal wb_in  : t_wishbone_master_in;
  signal wb_out : t_wishbone_master_out;

  signal irq_tx     : std_logic;
  signal irq_rx_ack : std_logic;
  signal irq_rx     : std_logic;

  signal nrx_newpacket, nrx_newpacket_d0 : std_logic;

  signal irq_txts    : std_logic;
  signal irq_tx_ack  : std_logic;
  signal irq_tx_mask : std_logic;

  signal txtsu_ack_int : std_logic;

begin  -- behavioral


-----------------------------------------------------------------------------
-- memory access arbitration
-----------------------------------------------------------------------------

  arbitrate_mem : process(clk_sys_i, rst_n_i)
  begin
    if rising_edge(clk_sys_i) then
      if rst_n_i = '0' then
        mem_arb_rx <= '0';
      else
        mem_arb_rx <= not mem_arb_rx;
      end if;
    end if;
  end process;

  mem_arb_tx <= not mem_arb_rx;
  mem_addr_o <= std_logic_vector(ntx_mem_a) when mem_arb_rx = '0' else std_logic_vector(nrx_mem_a);
  mem_data_o <= (others => '0')             when nrx_mux_d = '0'
                else nrx_mem_d;
  ntx_mem_d <= mem_data_i;
  mem_wr_o  <= nrx_mem_wr when mem_arb_rx = '1' else '0';

-------------------------------------------------------------------------------
-- TX Path  (Host -> Fabric)
-------------------------------------------------------------------------------  

-- helper signals to avoid big IF conditions in the FSM
  ntx_cntr_is_zero    <= '1' when (ntx_cntr = to_unsigned(0, ntx_cntr'length))       else '0';
  ntx_cntr_is_one     <= '1' when (ntx_cntr = to_unsigned(1, ntx_cntr'length))       else '0';
  ntx_ackcntr_is_zero <= '1' when (ntx_ackcntr = to_unsigned(0, ntx_ackcntr'length)) else '0';
  ntx_timeout_is_zero <= '1' when (ntx_timeout = to_unsigned(0, ntx_timeout'length)) else '0';

  tx_fsm : process(clk_sys_i, rst_n_i)
  begin
    if rising_edge(clk_sys_i) then
      if rst_n_i = '0' then
        src_dat_o          <= (others => '0');
        src_adr_o          <= (others => '0');
        src_cyc_o          <= '0';
        src_stb_o          <= '0';
        irq_tx             <= '0';
        ntx_has_oob        <= '0';
        ntx_mem_a          <= (others => '0');
        ntx_cntr           <= (others => '0');
        ntx_ackcntr        <= (others => '0');
        ntx_data_reg       <= (others => '0');
        ntx_status_reg     <= (others => '0');
        ntx_start_delayed  <= '0';
        ntx_state          <= TX_IDLE;

        regs_in.mcr_tx_error_i <= '0';
        regs_in.mcr_tx_idle_i  <= '0';

      else
        case ntx_state is

-------------------------------------------------------------------------------
-- Idle state: we wait until the host starts the DMA transfer
-------------------------------------------------------------------------------
          when TX_IDLE =>
            src_cyc_o <= '0';
            src_stb_o <= '0';
            -- keep the TX start bit (it's active for single clock cycle) in
            -- case we needed to align the FSM cycle with the memory arbiter
            if(regs_out.mcr_tx_start_o = '1') then
              ntx_start_delayed <= '1';
            end if;

            -- TX interrupt is disabled. Just assert the TX_IDLE.
            if(irq_tx_mask = '0') then
              regs_in.mcr_tx_idle <= '1';
            elsif(irq_tx_ack = '1') then
              irq_tx            <= '0';
              regs_in.mcr_tx_idle <= '1';
            end if;

            -- initialize timeout of TX_END_PACKET
            ntx_timeout <= to_unsigned(100, ntx_timeout'length);

            -- the host loaded new TX DMA buffer address
            if(regs_out.tx_addr_load = '1') then
              ntx_mem_a <= unsigned(regs_out.tx_addr_new(g_memsize_log2+1 downto 2));
            end if;

            -- the host started the DMA xfer (and we are "phased" with the arbiter)
            if(src_err_i = '0' and ntx_start_delayed = '1' and mem_arb_tx = '0') then
              ntx_state          <= TX_READ_DESC;
              -- clear the TX flags
              regs_in.mcr_tx_error <= '0';
              regs_in.mcr_tx_idle  <= '0';
            end if;


-------------------------------------------------------------------------------
-- Read descriptor header state: check if there's another descriptor in the buffer
-- and eventually, start transmitting it
-------------------------------------------------------------------------------
          when TX_READ_DESC =>
            ntx_start_delayed <= '0';

            if(mem_arb_tx = '0') then   -- memory is ready?
              -- feed the current TX DMA address as the readback value of TX_ADDR Wishbone
              -- register
              regs_in.tx_addr_cur(g_memsize_log2+1 downto 0)                      <= std_logic_vector(ntx_mem_a) & "00";
              regs_in.tx_addr_cur(regs_in.tx_addr_cur'high downto g_memsize_log2+2) <= (others => '0');

              -- if we have no more valid TX descriptors, trigger an interrupt and wait for
              -- another DMA transfer
              if(ntx_desc_valid = '0') then
                ntx_state <= TX_IDLE;
                irq_tx    <= '1';
              else
                -- read the descriptor contents (size, 802.1q/OOB enables)
                ntx_size_odd     <= ntx_desc_odd;
                ntx_cntr         <= unsigned(ntx_desc_size);
                ntx_ackcntr      <= unsigned(ntx_desc_size) + 1;  --+1 for status reg
                ntx_has_oob      <= ntx_desc_with_oob;
                ntx_status_hp    <= '0';
                ntx_status_smac  <= ntx_desc_has_src_mac;
                ntx_status_crc   <= '0';
                ntx_status_err   <= '0';
                ntx_status_class <= c_CLASS_PTP;
                ntx_state        <= TX_STATUS;
                ntx_mem_a        <= ntx_mem_a + 1;
              end if;
            end if;

-------------------------------------------------------------------------------
-- State status: send status word
-------------------------------------------------------------------------------
          when TX_STATUS =>

            src_cyc_o <= '1';
            src_stb_o <= '1';
            src_adr_o <= c_WBP_STATUS;
            if(src_stall_i = '0') then
              src_dat_o <= ntx_status_reg;
              ntx_state <= TX_START_PACKET;
            end if;

            if(src_ack_i = '1') then
              ntx_ackcntr <= ntx_ackcntr - 1;
            end if;

-------------------------------------------------------------------------------
-- Start packet state: asserts CYC signal and reads first word to transmit
-------------------------------------------------------------------------------            
          when TX_START_PACKET =>

            src_cyc_o <= '1';
            src_stb_o <= '0';
            -- check if the memory is ready, read the 1st word of the payload
            if(src_stall_i = '0' and mem_arb_tx = '0') then
              ntx_data_reg <= f_buf_swap_endian_32(ntx_mem_d);
              src_cyc_o    <= '1';
              ntx_state    <= TX_HWORD;
              ntx_mem_a    <= ntx_mem_a + 1;
            end if;


--------------------------------------------------------------------------------
-- State "Transmit HI word" - transmit the most significant word of the packet
-------------------------------------------------------------------------------
          when TX_HWORD =>
            ntx_curst <= TX_HWORD;

            src_cyc_o <= '1';
            src_stb_o <= '1';
            if(src_err_i = '1') then
              regs_in.mcr_tx_error <= '1';
              irq_tx             <= '1';
              ntx_state          <= TX_IDLE;
            end if;

            if(ntx_cntr_is_zero = '1' and ntx_has_oob = '1') then
              src_adr_o <= c_WBP_OOB;
            else
              src_adr_o <= c_WBP_DATA;
            end if;

            if(src_err_i = '0' and src_stall_i = '0') then
              src_dat_o <= ntx_data_reg(31 downto 16);
              if(ntx_cntr_is_zero = '1') then
                ntx_cntr  <= to_unsigned(c_GAP_SIZE, ntx_cntr'length);
                src_stb_o <= '0';
                ntx_state <= TX_END_PACKET;
              elsif(ntx_cntr = to_unsigned(1, ntx_cntr'length)) then
                --seems like odd number of words, so don't send here, prepare 
                --immediately new word and jump to TX_LWORD to send it out
                src_stb_o <= '0';
                if(ntx_has_oob = '1') then
                  src_adr_o <= c_WBP_OOB;
                end if;
                src_dat_o <= ntx_data_reg(15 downto 0);
                ntx_state <= TX_LWORD;
              else
                ntx_cntr  <= ntx_cntr - 1;
                ntx_state <= TX_LWORD;
              end if;
            end if;

            if(src_ack_i = '1') then
              ntx_ackcntr <= ntx_ackcntr - 1;
            end if;

--------------------------------------------------------------------------------
-- State "Transmit LO word" - transmit the least significant word of the packet
-------------------------------------------------------------------------------
          when TX_LWORD =>
            ntx_curst <= TX_LWORD;

            src_cyc_o <= '1';
            src_stb_o <= '1';
            src_stb_o <= '1';
            if(src_err_i = '1') then
              regs_in.mcr_tx_error <= '1';
              irq_tx             <= '1';
              ntx_state          <= TX_IDLE;
            end if;

            --set OOB adr when we are sending last word of the packet, descriptor says there is oob and
            --there was a immediate jump from TX_HWORD(odd number of words) or there is no stall
            --why? because if there was no immediate jump and STALL='1' then we have to remain with c_WBP_DATA
            --so that Slave could get the word sent by TX_HWORD after deactivating STALL
            if(ntx_cntr_is_one = '1' and ntx_has_oob = '1' and (ntx_size_odd = '1' or src_stall_i = '0')) then
              src_adr_o <= c_WBP_OOB;
            else
              src_adr_o <= c_WBP_DATA;
            end if;

            -- the TX fabric is ready, the memory is ready and we haven't reached the end
            -- of the packet yet:

            if(src_stall_i = '0') then
              src_dat_o <= ntx_data_reg (15 downto 0);
              if(mem_arb_tx = '0' and ntx_cntr_is_one = '0') then
                ntx_data_reg <= f_buf_swap_endian_32(ntx_mem_d);
                ntx_cntr     <= ntx_cntr - 1;
                ntx_mem_a    <= ntx_mem_a + 1;
                ntx_state    <= TX_HWORD;

              elsif(ntx_cntr_is_one = '1') then
                -- We're at the end of the packet
                ntx_cntr  <= to_unsigned(c_GAP_SIZE, ntx_cntr'length);
                src_stb_o <= '1';
                ntx_state <= TX_END_PACKET;
              else
                src_stb_o <= '0';
              end if;
            elsif(src_stall_i = '1' and ntx_cntr_is_one = '1' and ntx_size_odd = '1') then
              src_dat_o <= ntx_data_reg(15 downto 0);
              ntx_cntr  <= to_unsigned(c_GAP_SIZE, ntx_cntr'length);
              ntx_state <= TX_END_PACKET;
            else
              ntx_state <= TX_LWORD;
            end if;

            if(src_ack_i = '1') then
              ntx_ackcntr <= ntx_ackcntr - 1;
            end if;

-------------------------------------------------------------------------------
-- State end-of-packet: wait for ACKs and generate an inter-packet gap
-------------------------------------------------------------------------------
          when TX_END_PACKET =>
            ntx_curst <= TX_END_PACKET;

            src_stb_o <= '0';
            if(src_stall_i = '1' and ntx_ackcntr_is_zero = '0') then
              src_stb_o <= '1';
            else
              --inter-packet gap generation
              if(ntx_cntr_is_zero = '0') then
                ntx_cntr <= ntx_cntr - 1;
              end if;
              --ACKs reception
              if(src_ack_i = '1') then
                ntx_ackcntr <= ntx_ackcntr - 1;
              end if;
              --disable CYC if all ACKs received
              if(ntx_ackcntr_is_zero = '1') then
                src_cyc_o <= '0';
              end if;
              --timeout in case something went wrong and we won't ever
              --get those ACKs
              if(ntx_timeout_is_zero = '1') then
                regs_in.mcr_tx_error <= '1';
              else
                ntx_timeout <= ntx_timeout - 1;
              end if;
              --finish when gap generated and all ACKs received or timeout expired
              if(ntx_cntr_is_zero = '1' and (ntx_ackcntr_is_zero = '1' or minic_mcr_tx_error = '1')) then
                ntx_state <= TX_READ_DESC;
              end if;
            end if;
          when others => null;
        end case;
      end if;
    end if;
  end process;

-- these are never used:
  src_sel_o <= "11";
  src_we_o  <= '1';

-------------------------------------------------------------------------------
-- RX Path (Fabric ->  Host)
-------------------------------------------------------------------------------  

  rx_fsm : process(clk_sys_i, rst_n_i)
  begin
    if rising_edge(clk_sys_i) then
      if rst_n_i = '0' then
        nrx_state      <= RX_WAIT_SOF;
        nrx_mem_a      <= (others => '0');
        nrx_mem_d      <= (others => '0');
        nrx_mux_d      <= '0';
        nrx_mem_wr     <= '0';
        nrx_avail      <= (others => '0');
        nrx_status_reg <= (others => '0');
        nrx_oob_reg    <= (others => '0');
        nrx_toggle     <= '0';
        nrx_stall_mask <= '0';
        nrx_bytesel    <= '0';
        nrx_size       <= (others => '0');
        nrx_acksize    <= (others => '0');
        nrx_buf_full   <= '0';
        nrx_has_oob    <= '0';

        regs_in.rx_addr_cur  <= (others => '0');
        regs_in.mcr_rx_ready <= '0';
        regs_in.mcr_rx_full  <= '0';
        nrx_newpacket      <= '0';

        snk_ack_o <= '0';
      else
        -- Host can modify the RX DMA registers only when the DMA engine is disabled
        -- (MCR_RX_EN = 0)
        if(regs_out.mcr_rx_en = '0') then

          nrx_newpacket      <= '0';
          -- mask out the stall line on the fabric I/F, so the endpoint
          -- can cut the traffic using 802.1 flow control
          nrx_stall_mask     <= '0';
          nrx_state          <= RX_WAIT_SOF;
          regs_in.mcr_rx_ready <= '0';

          -- handle writes to RX_ADDR and RX_AVAIL
          if(regs_out.rx_addr_load = '1') then
            nrx_mem_a_saved   <= unsigned(minic_rx_addr_new(g_memsize_log2+1 downto 2));
            regs_in.rx_addr_cur <= (others => '0');
          end if;

          if(regs_out.rx_avail_load = '1') then
            nrx_buf_full      <= '0';
            regs_in.mcr_rx_full <= '0';
            nrx_avail         <= unsigned(regs_out.rx_avail_new(nrx_avail'high downto 0));
          end if;

          snk_ack_o <= '0';
        else

          case nrx_state is

-------------------------------------------------------------------------------
-- State "Wait for start of frame". We wait until CYC goes high
-- on the RX fabric and then we commence reception of the packet.
-------------------------------------------------------------------------------
            when RX_WAIT_SOF =>

              nrx_newpacket <= '0';
              nrx_mem_wr    <= '0';
              nrx_has_oob   <= '0';
              nrx_bytesel   <= '0';
              nrx_size      <= (others => '0');
              if(g_buffer_little_endian = false) then
                nrx_mem_d(15 downto 0) <= snk_dat_i;
              else
                nrx_mem_d(15 downto 8) <= snk_dat_i(7 downto 0);
                nrx_mem_d(7 downto 0)  <= snk_dat_i(15 downto 8);
              end if;
              nrx_mux_d   <= '0';
              nrx_mem_a   <= nrx_mem_a_saved;
              nrx_toggle  <= '0';
              snk_ack_o   <= '0';
              nrx_acksize <= (others => '0');

              regs_in.mcr_rx_full <= nrx_buf_full;

              if(snk_cyc_i = '1') then
                nrx_size       <= nrx_size + 1;
                nrx_stall_mask <= '0';
                nrx_state      <= RX_ALLOCATE_DESCRIPTOR;
              else
                nrx_stall_mask <= not nrx_buf_full;
              end if;

-------------------------------------------------------------------------------
-- State "Allocate RX descriptor": puts an empty (invalid) RX descriptor at the
-- current location in the RX buffer and then starts receiving the data
-------------------------------------------------------------------------------              
            when RX_ALLOCATE_DESCRIPTOR =>

              snk_ack_o  <= '0';
              nrx_toggle <= '1';

              -- wait until we have memory access
              if(mem_arb_rx = '0') then
                nrx_mem_a_saved <= nrx_mem_a;
                nrx_avail       <= nrx_avail - 1;
                nrx_mux_d       <= '0';
                nrx_mem_wr      <= '1';

                snk_ack_o   <= '1';
                nrx_acksize <= nrx_acksize + 1;

                nrx_state      <= RX_DATA;
                -- allow the fabric to receive the data
                nrx_stall_mask <= '1';
              end if;

-------------------------------------------------------------------------------
-- State "Receive data". Receive data, write it into the DMA memory
-------------------------------------------------------------------------------              
            when RX_DATA =>

              nrx_mux_d  <= '1';
              nrx_mem_wr <= '0';

              -- if we have no more space in memory then generate error
              -- and finish reception
              if(nrx_avail = to_unsigned(0, nrx_avail'length)) then
                nrx_status_err <= '1';
                nrx_buf_full   <= '1';
                nrx_state      <= RX_UPDATE_DESC;
              end if;

              -- error/end-of-frame?
              if(snk_cyc_i = '0' or nrx_status_err = '1') then
                snk_ack_o <= '0';

                -- flush the remaining packet data into the DMA buffer
                nrx_state <= RX_MEM_FLUSH;

                if(g_buffer_little_endian = false) then
                  if (nrx_toggle = '1') then
                    nrx_mem_a               <= nrx_mem_a + 1;
                    nrx_mem_d(31 downto 16) <= nrx_oob_reg;
                    nrx_mem_d(15 downto 0)  <= (others => '0');
                  else
                    nrx_mem_d(15 downto 0) <= nrx_oob_reg;
                  end if;
                else
                  if (nrx_toggle = '1') then
                    nrx_mem_d(31 downto 24) <= nrx_oob_reg(7 downto 0);
                    nrx_mem_d(23 downto 16) <= nrx_oob_reg(15 downto 8);
                  else
                    nrx_mem_a               <= nrx_mem_a + 1;
                    nrx_mem_d(31 downto 16) <= (others => '0');
                    nrx_mem_d(15 downto 8)  <= nrx_oob_reg(7 downto 0);
                    nrx_mem_d(7 downto 0)   <= nrx_oob_reg(15 downto 8);
                  end if;
                end if;

                -- disable the RX fabric reception, so we won't get another
                -- packet before we are done with the RX descriptor update
                nrx_stall_mask <= '0';
              end if;


              if(snk_stb_i = '1') then

                -- latch the bytesel signal to support frames having odd lengths
                if(snk_sel_i = "10") then
                  nrx_bytesel <= '1';
                end if;

                snk_ack_o   <= '1';
                nrx_acksize <= nrx_acksize + 1;

                --================--
                ----  DATA REG  ----
                if(snk_adr_i = c_WBP_DATA) then
                  nrx_size <= nrx_size + 1;
                  -- pack two 16-bit words received from the fabric I/F into one
                  -- 32-bit DMA memory word
                  if(g_buffer_little_endian = false) then
                    -- big endian RX buffer
                    if(nrx_toggle = '0') then
                      nrx_mem_d(31 downto 16) <= snk_dat_i;
                    else
                      nrx_mem_d(15 downto 0) <= snk_dat_i;
                    end if;
                  else
                    -- little endian RX buffer
                    if(nrx_toggle = '0') then
                      nrx_mem_d(15 downto 8) <= snk_dat_i(7 downto 0);
                      nrx_mem_d(7 downto 0)  <= snk_dat_i(15 downto 8);
                    else
                      nrx_mem_d(31 downto 24) <= snk_dat_i(7 downto 0);
                      nrx_mem_d(23 downto 16) <= snk_dat_i(15 downto 8);
                    end if;
                  end if;
                  nrx_toggle <= not nrx_toggle;
                --================--
                ---- STATUS REG ----
                elsif(snk_adr_i = c_WBP_STATUS) then
                  if(g_buffer_little_endian = false) then
                    nrx_status_reg(15 downto 8) <= snk_dat_i(7 downto 0);
                    nrx_status_reg(7 downto 0)  <= snk_dat_i(15 downto 8);
                  else
                    nrx_status_reg(15 downto 0) <= snk_dat_i(15 downto 0);
                  end if;
                --===============--
                ------- OOB -------
                elsif(snk_adr_i = c_WBP_OOB) then
                  nrx_size    <= nrx_size + 1;
                  -- we've got RX OOB tag? Remember it and later put it in the
                  -- descriptor header
                  nrx_has_oob <= '1';
                  if(g_buffer_little_endian = false) then
                    nrx_oob_reg(15 downto 8) <= snk_dat_i(7 downto 0);
                    nrx_oob_reg(7 downto 0)  <= snk_dat_i(15 downto 8);
                  else
                    nrx_oob_reg(15 downto 0) <= snk_dat_i(15 downto 0);
                  end if;
                end if;
              elsif(snk_stb_i = '0') then
                snk_ack_o <= '0';
              end if;

              -- we've got the second valid word of the payload, write it to the
              -- memory
              if(nrx_avail /= to_unsigned(0, nrx_avail'length) and nrx_toggle = '1' and snk_stb_i = '1' and snk_cyc_i = '1') then
                nrx_mem_a  <= nrx_mem_a + 1;
                nrx_mem_wr <= '1';
                nrx_avail  <= nrx_avail - 1;

                -- check if we are synchronized with the memory write arbiter.
                if(mem_arb_rx = '1') then
                  nrx_state <= RX_MEM_RESYNC;
                end if;
              else
                -- nothing to write
                nrx_mem_wr <= '0';
              end if;

-------------------------------------------------------------------------------
-- State "Memory resync": a "wait state" entered when the miNIC tries to write the RX
-- payload, but the memory access is given for the TX path at the moment.
-------------------------------------------------------------------------------
            when RX_MEM_RESYNC =>
              snk_ack_o <= '0';
              nrx_state <= RX_DATA;

-------------------------------------------------------------------------------
-- State "Memory flush": flushes the remaining contents of RX data register
-- into the DMA buffer after end-of-packet
-------------------------------------------------------------------------------
            when RX_MEM_FLUSH =>
              snk_ack_o  <= '0';
              nrx_mem_wr <= '1';
              if(mem_arb_rx = '0') then
                nrx_avail <= nrx_avail - 1;
                nrx_state <= RX_UPDATE_DESC;
              end if;

-------------------------------------------------------------------------------
-- State "Update RX descriptor": writes the frame size, OOB presence and error
-- flags into the empty RX descriptor allocated at the beginning of the reception
-- of the frame, and marks the descriptor as valid. Also triggers the RX ready
-- interrupt.
-------------------------------------------------------------------------------
              
            when RX_UPDATE_DESC =>
              snk_ack_o <= '0';

              ------------------------------------
              -- Discard packets other than PTP --
              ------------------------------------
              if(nrx_status_class /= c_CLASS_PTP) then
                nrx_mem_wr         <= '0';
                nrx_newpacket      <= '0';
                regs_in.mcr_rx_ready <= '0';
                nrx_state          <= RX_WAIT_SOF;
              elsif(mem_arb_rx = '0') then

                -- store the current write pointer as a readback value of RX_ADDR register, so
                -- the host can determine the RX descriptor we're actually working on
                regs_in.rx_addr_cur(g_memsize_log2+1 downto 0)                      <= std_logic_vector(nrx_mem_a_saved) & "00";
                regs_in.rx_addr_cur(regs_in.rx_addr_cur'high downto g_memsize_log2+2) <= (others => '0');

                nrx_mem_a       <= nrx_mem_a_saved;
                nrx_mem_a_saved <= nrx_mem_a + 1;

                -- compose the RX descriptor
                nrx_mem_d(31)                         <= '1';
                nrx_mem_d(30)                         <= nrx_status_err;
                nrx_mem_d(29)                         <= nrx_has_oob;
                nrx_mem_d(28 downto g_memsize_log2+1) <= (others => '0');
                nrx_mem_d(g_memsize_log2 downto 1)    <= std_logic_vector(nrx_size);
                nrx_mem_d(0)                          <= nrx_bytesel;

                nrx_mem_wr <= '1';

                -- trigger the RX interrupt and assert RX_READY flag to inform
                -- the host that we've received something
                nrx_newpacket      <= '1';
                regs_in.mcr_rx_ready <= '1';

                -- wait for another packet
                nrx_state <= RX_WAIT_SOF;
              else
                nrx_mem_wr <= '0';
              end if;
              
            when others => null;
          end case;
        end if;
      end if;
    end if;
  end process;

  snk_err_o <= nrx_buf_full;

-------------------------------------------------------------------------------
-- helper process for producing the RX fabric data request signal (combinatorial)
-------------------------------------------------------------------------------  
  gen_rx_dreq : process(nrx_stall_mask, nrx_state, mem_arb_rx, nrx_toggle, regs_out.mcr_rx_en)
  begin
    -- make sure we don't have any incoming data when the reception is masked (e.g.
    -- the miNIC is updating the descriptors of finishing the memory write. 
    if(regs_out.mcr_rx_en = '0' or nrx_state = RX_ALLOCATE_DESCRIPTOR or nrx_state = RX_UPDATE_DESC or nrx_state = RX_MEM_FLUSH) then
      snk_stall_o <= '1';
    elsif(nrx_stall_mask = '0') then
      snk_stall_o <= '0';

    -- the condition below forces the RX FSM to go into RX_MEM_RESYNC state. Don't
    -- receive anything during this time
    elsif(nrx_toggle = '1' and mem_arb_rx = '1') then
      snk_stall_o <= '1';
    else
      snk_stall_o <= '0';
    end if;
  end process;


-------------------------------------------------------------------------------
-- TX Timestamping unit
-------------------------------------------------------------------------------  
  tsu_fsm : process(clk_sys_i, rst_n_i)
  begin
    if rising_edge(clk_sys_i) then
      if(rst_n_i = '0') then
        minic_tsfifo_wr_req <= '0';
        minic_tsfifo_fid    <= (others => '0');
        minic_tsfifo_pid    <= (others => '0');
        minic_tsfifo_tsval  <= (others => '0');
        txtsu_ack_int       <= '0';
      else
        -- Make sure the timestamp is written to the FIFO only once.

        if(txtsu_valid_i = '1' and txtsu_ack_int = '0' and minic_tsfifo_wr_full = '0') then
          minic_tsfifo_wr_req <= '1';
          minic_tsfifo_tsval  <= txtsu_tsval_i;
          minic_tsfifo_fid    <= txtsu_frame_id_i;
          minic_tsfifo_pid    <= txtsu_port_id_i;
          txtsu_ack_int       <= '1';
        else
          txtsu_ack_int       <= '0';
          minic_tsfifo_wr_req <= '0';
        end if;
      end if;
    end if;
  end process;

  txtsu_ack_o <= txtsu_ack_int;

  handle_rx_interrupt : process(clk_sys_i, rst_n_i)
  begin
    if rising_edge(clk_sys_i) then
      if rst_n_i = '0' then
        irq_rx           <= '0';
        nrx_newpacket_d0 <= '0';
      else
        nrx_newpacket_d0 <= nrx_newpacket;

        if (nrx_newpacket_d0 = '0' and nrx_newpacket = '1') then
          irq_rx <= '1';
        elsif (regs_out.mcr_rx_full = '1') then
          irq_rx <= '1';
        elsif (irq_rx_ack = '1') then
          irq_rx <= '0';
        end if;
      end if;
    end if;
  end process;

  irq_txts <= not minic_tsfifo_wr_empty;


  U_Slave_Adapter : wb_slave_adapter
    generic map (
      g_master_use_struct  => true,
      g_master_mode        => CLASSIC,
      g_master_granularity => WORD,
      g_slave_use_struct   => false,
      g_slave_mode         => g_interface_mode,
      g_slave_granularity  => g_address_granularity)
    port map (
      clk_sys_i  => clk_sys_i,
      rst_n_i    => rst_n_i,
      sl_adr_i   => wb_adr_i,
      sl_dat_i   => wb_dat_i,
      sl_sel_i   => wb_sel_i,
      sl_cyc_i   => wb_cyc_i,
      sl_stb_i   => wb_stb_i,
      sl_we_i    => wb_we_i,
      sl_dat_o   => wb_dat_o,
      sl_ack_o   => wb_ack_o,
      sl_stall_o => wb_stall_o,
      master_i   => wb_in,
      master_o   => wb_out);

  U_WB_Slave : minic_wb_slave
    port map (
      rst_n_i          => rst_n_i,
      wb_clk_i         => clk_sys_i,
      wb_addr_i        => wb_out.adr(3 downto 0),
      wb_data_i        => wb_out.dat,
      wb_data_o        => wb_in.dat,
      wb_cyc_i         => wb_out.cyc,
      wb_sel_i         => wb_out.sel,
      wb_stb_i         => wb_out.stb,
      wb_we_i          => wb_out.we,
      wb_ack_o         => wb_in.ack,
      wb_irq_o         => wb_irq_o,
      tx_ts_read_ack_o => open,
      irq_tx_i         => irq_tx,
      irq_tx_ack_o     => irq_tx_ack,
      irq_tx_mask_o    => irq_tx_mask,
      irq_rx_i         => irq_rx,
      irq_rx_ack_o     => irq_rx_ack,
      irq_txts_i       => irq_txts);


  minic_rx_avail_cur (nrx_avail'high downto 0)                         <= std_logic_vector(nrx_avail);
  minic_rx_avail_cur (minic_rx_avail_cur'high downto nrx_avail'high+1) <= (others => '0');

end behavioral;
